----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    02:42:27 10/18/2021 
-- Design Name: 
-- Module Name:    task_1_bex_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity task_1_bex_1 is
    Port ( Q : out  STD_LOGIC;
           nQ : out  STD_LOGIC);
end task_1_bex_1;

architecture Behavioral of task_1_bex_1 is

signal a, b: std_logic;

begin

	a <= not b;
	b <= not a;
	
	nQ <= a;
	Q <= b;

end Behavioral;

